module cache_controller (
    input logic clk,
    input rst,
    input logic req_valid,
    input logic req_type,          // 0 = Read, 1 = Write
    input logic hit,
    input logic dirty_bit,
    input logic ready_mem,
    input logic acknowledge,
    output logic read_en_mem,
    output logic write_en_mem,
    output logic write_en,
    output logic read_en_cache,
    output logic refill,
    output logic done_cache
);

    typedef enum logic [2:0] {
        IDLE,
        COMPARE,
        WRITE_BACK,
        WRITE_ALLOCATE
    } state_t;

    state_t current_state, next_state;

    // State register
    always @(posedge clk or posedge rst) begin
        if (rst)
            current_state <= IDLE;
        else
            current_state <= next_state;
    end

    // Mealy outputs and state transitions
    always @(*) begin
        // Default values (safe defaults)
        read_en_mem    = 0;
        write_en_mem   = 0;
        write_en       = 0;
        read_en_cache  = 0;
        refill         = 0;
        acknowledge    = 0;
        next_state     = current_state;

        case (current_state)
            IDLE: begin
                if (req_valid)
                    next_state = COMPARE;
            end

            COMPARE: begin
                if (req_type == 0 && hit) begin
                    read_en_cache = 1;
                    done_cache = 1;
                    next_state = IDLE;
                end
                else if (req_type == 0 && !hit && dirty_bit) begin
                    write_en_mem = 1;            // Write dirty block to main memory
                    next_state = WRITE_BACK;
                end
                else if (req_type == 0 && !hit && !dirty_bit) begin
                    read_en_mem = 1;
                    next_state = WRITE_ALLOCATE;
                end
                else if (req_type == 1 && hit) begin
                    write_en = 1;  // allow CPU to write into cache
                    done_cache = 1;
                    next_state = IDLE;
                end
                else if (req_type == 1 && !hit && dirty_bit) begin
                    write_en_mem = 1;
                    next_state = WRITE_BACK;
                end
                else if (req_type == 1 && !hit && !dirty_bit) begin
                    read_en_mem = 1;
                    next_state = WRITE_ALLOCATE;
                end
            end

            WRITE_BACK: begin
                if (acknowledge) begin
                    read_en_mem = 1;
                    next_state = WRITE_ALLOCATE;
                end
            end

            WRITE_ALLOCATE: begin
                if (ready_mem) begin
                    refill = 1;
                    if (req_type == 0)
                        read_en_cache = 1;
                    else if (req_type == 1)
                        write_en = 1;
                    done_cache = 1;
                    next_state = IDLE;
                end
            end

            default: next_state = IDLE;
        endcase
    end

endmodule
